`timescale 1ns / 1ps

module IDU_tb;

	// Inputs
	reg [31:0] IR;

	// Outputs
	wire [7:0] IRN;
	wire [3:0] IRType;
	wire Unknown;

	// Instantiate the Unit Under Test (UUT)
	IDU uut (
		.IR(IR), 
		.IRN(IRN), 
		.IRType(IRType), 
		.Unknown(Unknown)
	);

	initial begin
		// Initialize Inputs
		IR = 0;

		IR = 32'h00430820;
		#10;
		IR = 32'h00430821;
		#10;
		IR = 32'h00430822;
		#10;
		IR = 32'h00430823;
		#10;
		IR = 32'h00020800;
		#10;
		IR = 32'h00020802;
		#10;
		IR = 32'h00020803;
		#10;
		IR = 32'h00620804;
		#10;
		IR = 32'h00620806;
		#10;
		IR = 32'h00620807;
		#10;
		IR = 32'h00430824;
		#10;
		IR = 32'h00430825;
		#10;
		IR = 32'h00430826;
		#10;
		IR = 32'h00430827;
		#10;
		IR = 32'h0043082a;
		#10;
		IR = 32'h0043082b;
		#10;
		IR = 32'h00220018;
		#10;
		IR = 32'h00220019;
		#10;
		IR = 32'h0022001a;
		#10;
		IR = 32'h0022001b;
		#10;
		IR = 32'h00200011;
		#10;
		IR = 32'h00200013;
		#10;
		IR = 32'h00000810;
		#10;
		IR = 32'h00000812;
		#10;
		IR = 32'h20410000;
		#10;
		IR = 32'h24410000;
		#10;
		IR = 32'h30410000;
		#10;
		IR = 32'h34410000;
		#10;
		IR = 32'h38410000;
		#10;
		IR = 32'h3c010000;
		#10;
		IR = 32'h28410000;
		#10;
		IR = 32'h2c410000;
		#10;
		IR = 32'h8c410000;
		#10;
		IR = 32'h80410000;
		#10;
		IR = 32'h90410000;
		#10;
		IR = 32'h84410000;
		#10;
		IR = 32'h94410000;
		#10;
		IR = 32'hac410000;
		#10;
		IR = 32'ha4410000;
		#10;
		IR = 32'ha0410000;
		#10;
		IR = 32'h10220009;
		#10;
		IR = 32'h14220008;
		#10;
		IR = 32'h18200007;
		#10;
		IR = 32'h1c200006;
		#10;
		IR = 32'h04200005;
		#10;
		IR = 32'h04210004;
		#10;
		IR = 32'h08000c32;
		#10;
		IR = 32'h0c000c32;
		#10;
		IR = 32'h03e00008;
		#10;
		IR = 32'h00400809;
		#10;
        
		// Add stimulus here

	end
      
endmodule

